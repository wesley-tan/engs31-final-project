-------------------------------------------------------------------------------
--  tb_top_morse.vhd
-------------------------------------------------------------------------------
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity tb_top_morse is
end entity;

architecture sim of tb_top_morse is

  -----------------------------------------------------------------------------
  --  DUT component declaration
  -----------------------------------------------------------------------------
  component Top_Morse is
    port (
      clk       : in  std_logic;
      rx        : in  std_logic;
      led_out   : out std_logic;
      sound_out : out std_logic
    );
  end component;

  -----------------------------------------------------------------------------
  --  Simulation constants
  -----------------------------------------------------------------------------
  constant CLK_PERIOD  : time := 10 ns;           -- 1 MHz
  constant clk_period_divided : time := 1000 ns;
  constant BAUD_PERIOD: integer:= 104;      -- 9600 baud
    

  -----------------------------------------------------------------------------
  --  DUT I/O signals
  -----------------------------------------------------------------------------
  signal clk       : std_logic := '0';
  signal rx        : std_logic := '1';  -- UART line idles high
  signal led_out_s   : std_logic;
  signal sound_out_s : std_logic;

begin
  ---------------------------------------------------------------------------
  --  clock generator
  ---------------------------------------------------------------------------
   clk_process :process
    begin
        clk <= '0';
        wait for clk_period/2;
        clk <= '1';
        wait for clk_period/2;
    end process;

  ---------------------------------------------------------------------------
  --  DUT instantiation
  ---------------------------------------------------------------------------
  uut : Top_Morse
    port map (
      clk       => clk,
      rx        => rx,
      led_out   => led_out_s,
      sound_out => sound_out_s
    );

  ---------------------------------------------------------------------------
  --  Stimulus process : sends "SOS" over UART
  ---------------------------------------------------------------------------
  stim : process
    -------------------------------------------------------------------------
    -- helper to transmit one 8-N-1 UART byte (LSB first)
    -------------------------------------------------------------------------
   
    begin
    
             Rx <= '1';
        
        wait for clk_period_divided * 10;
        
        -- Scenario 1: Load data 
        Rx <= '0';  -- Load the data
        wait for BAUD_PERIOD* clk_period_divided;
        
        -- Scenario 2: Load data "11001100"
        Rx <= '1';  -- Load the data
        wait for BAUD_PERIOD* clk_period_divided;
        
        -- Scenario 2: Load data "11001100"
        Rx <= '0';  -- Load the data
        wait for BAUD_PERIOD* clk_period_divided;

        
        
                -- Scenario 2: Load data "11001100"
        Rx <= '0';  -- Load the data
        wait for BAUD_PERIOD* clk_period_divided;

        Rx <= '0';  -- Load the data
        wait for BAUD_PERIOD* clk_period_divided;
        
        Rx <= '1';  -- Load the data
        wait for BAUD_PERIOD* clk_period_divided;
        
        Rx <= '1';  -- Load the data  
        wait for BAUD_PERIOD* clk_period_divided;


        Rx <= '0';  -- Load the data
        wait for BAUD_PERIOD*clk_period_divided;
        
        Rx <= '0';  -- Load the data
        wait for BAUD_PERIOD*clk_period_divided;
        Rx <= '1';  -- Load the data
		wait for 2*BAUD_PERIOD*clk_period_divided;

        -- Restart Transmission
        Rx <= '0';  -- Load the data
        wait for BAUD_PERIOD* clk_period_divided;
        
        -- Scenario 2: Load data "11001100"
        Rx <= '1';  -- Load the data
        wait for BAUD_PERIOD* clk_period_divided;
        
        -- Scenario 2: Load data "11001100"
        Rx <= '1';  -- Load the data
        wait for BAUD_PERIOD* clk_period_divided;

        
        
                -- Scenario 2: Load data "11001100"
        Rx <= '1';  -- Load the data
        wait for BAUD_PERIOD* clk_period;

        Rx <= '0';  -- Load the data
        wait for BAUD_PERIOD* clk_period;
        
        Rx <= '1';  -- Load the data
        wait for BAUD_PERIOD* clk_period;
        
        Rx <= '0';  -- Load the data  
        wait for BAUD_PERIOD* clk_period;


        Rx <= '1';  -- Load the data
        wait for BAUD_PERIOD*clk_period;
        
        Rx <= '0';  -- Load the data
        wait for BAUD_PERIOD*clk_period;
        Rx <= '1';  -- Load the data
		
        
        wait;
 
  end process;

end architecture sim;
